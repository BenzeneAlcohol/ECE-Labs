module hmlo(A,B,C);
input A,B;
output C;
endmodule;